module top(
    input sysclk_n,
    input sysclk_p,
    output  :qw

